* G:\STUDY\CSE209\Project final Cse209.sch

* Schematics Version 9.1 - Web Update 1
* Thu Sep 09 11:01:15 2021


.PARAM         RVAR=10 

** Analysis setup **
.DC LIN PARAM RVAR 0.001 3.5 0.001 
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Project final Cse209.net"
.INC "Project final Cse209.als"


.probe


.END
